module for a 2-bit adder with carry-in and carry-out.

Inputs:
- a (1 bit)
- b (1 bit)
- cin (1 bit, carry-in)

Outputs:
- sum (1 bit)
- cout (1 bit, carry-out)

The module should be written in Verilog syntax:
module adder(
  input a,
  input b,
  input cin,
  output sum,
  output cout
);

endmodule