module that implements a 2-to-1 multiplexer.

Module requirements:
1. Inputs: a (1 bit), b (1 bit), sel (1 bit selector)
2. Output: y (1 bit output)

Use standard Verilog syntax and include 'assign' statement for logic.
Ensure the module starts with 'module' and ends with 'endmodule